/***************************************************
Student Name: 
Student ID: 
***************************************************/

`timescale 1ns/1ps

module Adder(
    input  [31:0] src1_i,
	input  [31:0] src2_i,
	output [31:0] sum_o
	);
    
/* Write your code HERE */



endmodule